`timescale 1ns/100ps

module halfadder(output s, output c, input a, input b);
	
